
module tb;
    hello dut ();

    initial begin
        $display ("hello TB 0-r1");
    end;

endmodule
