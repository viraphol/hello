
module tb;
    hello dut ();

    initial begin
        $display ("hello TB git-r1");
    end;

endmodule
