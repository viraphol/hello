
module tb_erupt;
    hello dut ();

    initial begin
        $display ("hello TB git-r1 erupt test");
    end;

endmodule
